library ieee;
use ieee.std_logic_1164.all;

entity my_entity is
port(
     port_name_1 : in std_logic   ;
     port_name2:   out std_logic  ;
     port_name3:   inout std_logic) ;

end my_entity;


     
