----Exercise 3.6----

library ieee;
use ieee.std_logic_1164.all;

entity sys1 is 
    port  (a_in1, b_in2, clk, ctrl_int: in  std_logic;
          out_b: out std_logic);

end sys1;

